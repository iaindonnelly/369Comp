`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11/08/2017 07:18:01 PM
// Design Name: 
// Module Name: top
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module top(Clk,Reset,Something);

input Clk,Reset;

output reg Something;
    wire  A1,B1,1Out;
    wire  A2,B2,2Out;
    wire  A3,B3,3Out;
    wire  A4,B4,4Out;
    wire  A5,B5,5Out;
    wire  A6,B6,6Out;
    wire  A7,B7,7Out;
    wire  A8,B8,8Out;
    wire  A9,B9,9Out;






    Sadder Sadder1(A1,B1,1Out);
    Sadder Sadder2(A2,B2,2Out);
    Sadder Sadder3(A3,B3,3Out);
    Sadder Sadder4(A4,B4,4Out);
    Sadder Sadder5(A5,B5,5Out);
    Sadder Sadder6(A6,B6,6Out);
    Sadder Sadder7(A7,B7,7Out);
    Sadder Sadder8(A8,B8,8Out);
    Sadder Sadder9(A9,B9,9Out);
    Sadder Sadder10(10A,10B,10Out);
    Sadder Sadder11(11A,11B,11Out);
    Sadder Sadder12(12A,12B,12Out);
    Sadder Sadder13(13A,13B,13Out);
    Sadder Sadder14(14A,14B,14Out);
    Sadder Sadder15(15A,15B,15Out);
    Sadder Sadder16(16A,16B,16Out);
    
    adder adder1(A,B,Out);
    adder adder2(A,B,Out);
    adder adder3(A,B,Out);
    adder adder4(A,B,Out);
    adder adder5(A,B,Out);
    adder adder6(A,B,Out);
    adder adder7(A,B,Out);
    adder adder8(A,B,Out);
    
    adder adder9(A,B,Out);
    adder adder10(A,B,Out);
    adder adder11(A,B,Out);
    adder adder12(A,B,Out);
    
    adder adder13(A,B,Out);
    adder adder14(A,B,Out);
    
    adder adder15(A,B,Out);


always@(*) begin 

end
endmodule
